

module tb;

    // Input
    reg [7:0] X;
    // Outputs
    wire [4:0] ones;
    CountOnes uut (
        .X(X), 
        .ones(ones)
    );

    initial begin
        X = 'b00000000;   #50;
        X = 'b00000001;   #50;
        X = 'b00000010;   #50;
        X = 'b00000011;   #50;
        X = 'b00000100;   #50;
        X = 'b00000101;   #50;
        X = 'b00000110;   #50;   
	X = 'b00000111;   #50;

	X = 'b00001000;   #50;
        X = 'b00001001;   #50;
        X = 'b00001010;   #50;
        X = 'b00001011;   #50;
        X = 'b00001100;   #50;
        X = 'b00001101;   #50;
        X = 'b00001110;   #50;   
	X = 'b00001111;   #50;

	X = 'b00010000;   #50;
        X = 'b00010001;   #50;
        X = 'b00010010;   #50;
        X = 'b00010011;   #50;
        X = 'b00010100;   #50;
        X = 'b00010101;   #50;
        X = 'b00010110;   #50;   
	X = 'b00010111;   #50;

	X = 'b00011000;   #50;
        X = 'b00011001;   #50;
        X = 'b00011010;   #50;
        X = 'b00011011;   #50;
        X = 'b00011100;   #50;
        X = 'b00011101;   #50;
        X = 'b00011110;   #50;   
	X = 'b00011111;   #50;

	X = 'b00100000;   #50;
        X = 'b00100001;   #50;
        X = 'b00100010;   #50;
        X = 'b00100011;   #50;
        X = 'b00100100;   #50;
        X = 'b00100101;   #50;
        X = 'b00100110;   #50;   
	X = 'b00100111;   #50;

	X = 'b00101000;   #50;
        X = 'b00101001;   #50;
        X = 'b00101010;   #50;
        X = 'b00101011;   #50;
        X = 'b00101100;   #50;
        X = 'b00101101;   #50;
        X = 'b00101110;   #50;   
	X = 'b00101111;   #50;

	X = 'b00110000;   #50;
        X = 'b00110001;   #50;
        X = 'b00110010;   #50;
        X = 'b00110011;   #50;
        X = 'b00110100;   #50;
        X = 'b00110101;   #50;
        X = 'b00110110;   #50;   
	X = 'b00110111;   #50;

	X = 'b00111000;   #50;
        X = 'b00111001;   #50;
        X = 'b00111010;   #50;
        X = 'b00111011;   #50;
        X = 'b00111100;   #50;
        X = 'b00111101;   #50;
        X = 'b00111110;   #50;   
	X = 'b00111111;   #50;

        X = 'b01000000;   #50;
        X = 'b01000001;   #50;
        X = 'b01000010;   #50;
        X = 'b01000011;   #50;
        X = 'b01000100;   #50;
        X = 'b01000101;   #50;
        X = 'b01000110;   #50;   
	X = 'b01000111;   #50;

	X = 'b01001000;   #50;
        X = 'b01001001;   #50;
        X = 'b01001010;   #50;
        X = 'b01001011;   #50;
        X = 'b01001100;   #50;
        X = 'b01001101;   #50;
        X = 'b01001110;   #50;   
	X = 'b01001111;   #50;

	X = 'b01010000;   #50;
        X = 'b01010001;   #50;
        X = 'b01010010;   #50;
        X = 'b01010011;   #50;
        X = 'b01010100;   #50;
        X = 'b01010101;   #50;
        X = 'b01010110;   #50;   
	X = 'b01010111;   #50;

	X = 'b01011000;   #50;
        X = 'b01011001;   #50;
        X = 'b01011010;   #50;
        X = 'b01011011;   #50;
        X = 'b01011100;   #50;
        X = 'b01011101;   #50;
        X = 'b01011110;   #50;   
	X = 'b01011111;   #50;

	X = 'b01100000;   #50;
        X = 'b01100001;   #50;
        X = 'b01100010;   #50;
        X = 'b01100011;   #50;
        X = 'b01100100;   #50;
        X = 'b01100101;   #50;
        X = 'b01100110;   #50;   
	X = 'b01100111;   #50;

	X = 'b01101000;   #50;
        X = 'b01101001;   #50;
        X = 'b01101010;   #50;
        X = 'b01101011;   #50;
        X = 'b01101100;   #50;
        X = 'b01101101;   #50;
        X = 'b01101110;   #50;   
	X = 'b01101111;   #50;

	X = 'b01110000;   #50;
        X = 'b01110001;   #50;
        X = 'b01110010;   #50;
        X = 'b01110011;   #50;
        X = 'b01110100;   #50;
        X = 'b01110101;   #50;
        X = 'b01110110;   #50;   
	X = 'b01110111;   #50;

	X = 'b01111000;   #50;
        X = 'b01111001;   #50;
        X = 'b01111010;   #50;
        X = 'b01111011;   #50;
        X = 'b01111100;   #50;
        X = 'b01111101;   #50;
        X = 'b01111110;   #50;   
	X = 'b01111111;   #50;

        X = 'b10000000;   #50;
        X = 'b10000001;   #50;
        X = 'b10000010;   #50;
        X = 'b10000011;   #50;
        X = 'b10000100;   #50;
        X = 'b10000101;   #50;
        X = 'b10000110;   #50;   
	X = 'b10000111;   #50;

	X = 'b10001000;   #50;
        X = 'b10001001;   #50;
        X = 'b10001010;   #50;
        X = 'b10001011;   #50;
        X = 'b10001100;   #50;
        X = 'b10001101;   #50;
        X = 'b10001110;   #50;   
	X = 'b10001111;   #50;

	X = 'b10010000;   #50;
        X = 'b10010001;   #50;
        X = 'b10010010;   #50;
        X = 'b10010011;   #50;
        X = 'b10010100;   #50;
        X = 'b10010101;   #50;
        X = 'b10010110;   #50;   
	X = 'b10010111;   #50;

	X = 'b10011000;   #50;
        X = 'b10011001;   #50;
        X = 'b10011010;   #50;
        X = 'b10011011;   #50;
        X = 'b10011100;   #50;
        X = 'b10011101;   #50;
        X = 'b10011110;   #50;   
	X = 'b10011111;   #50;

	X = 'b10100000;   #50;
        X = 'b10100001;   #50;
        X = 'b10100010;   #50;
        X = 'b10100011;   #50;
        X = 'b10100100;   #50;
        X = 'b10100101;   #50;
        X = 'b10100110;   #50;   
	X = 'b10100111;   #50;

	X = 'b10101000;   #50;
        X = 'b10101001;   #50;
        X = 'b10101010;   #50;
        X = 'b10101011;   #50;
        X = 'b10101100;   #50;
        X = 'b10101101;   #50;
        X = 'b10101110;   #50;   
	X = 'b10101111;   #50;

	X = 'b10110000;   #50;
        X = 'b10110001;   #50;
        X = 'b10110010;   #50;
        X = 'b10110011;   #50;
        X = 'b10110100;   #50;
        X = 'b10110101;   #50;
        X = 'b10110110;   #50;   
	X = 'b10110111;   #50;

	X = 'b10111000;   #50;
        X = 'b10111001;   #50;
        X = 'b10111010;   #50;
        X = 'b10111011;   #50;
        X = 'b10111100;   #50;
        X = 'b10111101;   #50;
        X = 'b10111110;   #50;   
	X = 'b10111111;   #50;

        X = 'b11000000;   #50;
        X = 'b11000001;   #50;
        X = 'b11000010;   #50;
        X = 'b11000011;   #50;
        X = 'b11000100;   #50;
        X = 'b11000101;   #50;
        X = 'b11000110;   #50;   
	X = 'b11000111;   #50;

	X = 'b11001000;   #50;
        X = 'b11001001;   #50;
        X = 'b11001010;   #50;
        X = 'b11001011;   #50;
        X = 'b11001100;   #50;
        X = 'b11001101;   #50;
        X = 'b11001110;   #50;   
	X = 'b11001111;   #50;

	X = 'b11010000;   #50;
        X = 'b11010001;   #50;
        X = 'b11010010;   #50;
        X = 'b11010011;   #50;
        X = 'b11010100;   #50;
        X = 'b11010101;   #50;
        X = 'b11010110;   #50;   
	X = 'b11010111;   #50;

	X = 'b11011000;   #50;
        X = 'b11011001;   #50;
        X = 'b11011010;   #50;
        X = 'b11011011;   #50;
        X = 'b11011100;   #50;
        X = 'b11011101;   #50;
        X = 'b11011110;   #50;   
	X = 'b11011111;   #50;

	X = 'b11100000;   #50;
        X = 'b11100001;   #50;
        X = 'b11100010;   #50;
        X = 'b11100011;   #50;
        X = 'b11100100;   #50;
        X = 'b11100101;   #50;
        X = 'b11100110;   #50;   
	X = 'b11100111;   #50;

	X = 'b11101000;   #50;
        X = 'b11101001;   #50;
        X = 'b11101010;   #50;
        X = 'b11101011;   #50;
        X = 'b11101100;   #50;
        X = 'b11101101;   #50;
        X = 'b11101110;   #50;   
	X = 'b11101111;   #50;

	X = 'b11110000;   #50;
        X = 'b11110001;   #50;
        X = 'b11110010;   #50;
        X = 'b11110011;   #50;
        X = 'b11110100;   #50;
        X = 'b11110101;   #50;
        X = 'b11110110;   #50;   
	X = 'b11110111;   #50;

	X = 'b11111000;   #50;
        X = 'b11111001;   #50;
        X = 'b11111010;   #50;
        X = 'b11111011;   #50;
        X = 'b11111100;   #50;
        X = 'b11111101;   #50;
        X = 'b11111110;   #50;   
	X = 'b11111111;   #50;


	

    end
      
endmodule